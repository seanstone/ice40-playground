module setbit(
  output LED1,
  output LED2,
  output LED3,
  output LED4,
  output LED5,
  output LED6,
  output LED7,
  output LED8
);

    wire LED1;
    wire LED2;
    wire LED3;
    wire LED4;
    wire LED5;
    wire LED6;
    wire LED7;
    wire LED8;

    assign LED1 = 1;
    assign LED2 = 0;
    assign LED3 = 0;
    assign LED4 = 0;
    assign LED5 = 0;
    assign LED6 = 0;
    assign LED7 = 0;
    assign LED8 = 0;

endmodule